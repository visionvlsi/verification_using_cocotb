`timescale 1ns / 1ps
module ary_mul(a,b,out);
input [7:0]a,b;
output [15:0]out;
wire c0,c1,c2,c3,c4,c5,c6,c7,c8,c9,c10,c11,c12,c13,c14,c15,c16,c17,c18,c19,c20,c21,c22,c23,c24,c25,c26,c27,c28,c29,c30,c31,c32,c33,c34,c35,c36,c37,c38,c39,c40,
c41,c42,c43,c44,c45,c46,c47,c48,c49,c50,c51,c52,c53,c54;
wire q1,q2,q3,q4,q5,q6,q7,q8,q9,q10,q11,q12,q13,q14,q15,q16,q17,q18,q19,q20,q21,q22,q23,q24,q25,q26,q27,q28,q29,q30,
     q31,q32,q33,q34,q35,q36,q37,q38,q39,q40,q41,q42,q43,q44,q45,q46,q47,q48,q49,q50,q51,q52,q53,q54,q55,q56,q57,q58,q59,q60,q61,q62,q63;
wire p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15;
wire s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,s13,s14,s15,s16,s17,s18,s19,s20,s21,s22,s23,s24,s25,s26,s27,s28,s29,s30,
     s31,s32,s33,s34,s35,s36,s37,s38,s39,s40,s41,s42;
	  
assign p0=a[0]&b[0],
		q1=a[0]&b[1],q2=a[0]&b[2],q3=a[0]&b[3],q4=a[0]&b[4],q5=a[0]&b[5],q6=a[0]&b[6],q7=a[0]&b[7],
		q8=a[1]&b[0],q9=a[1]&b[1],q10=a[1]&b[2],q11=a[1]&b[3],q12=a[1]&b[4],q13=a[1]&b[5],q14=a[1]&b[6],q15=a[1]&b[7],
		q16=a[2]&b[0],q17=a[2]&b[1],q18=a[2]&b[2],q19=a[2]&b[3],q20=a[2]&b[4],q21=a[2]&b[5],q22=a[2]&b[6],q23=a[2]&b[7],
		q24=a[3]&b[0],q25=a[3]&b[1],q26=a[3]&b[2],q27=a[3]&b[3],q28=a[3]&b[4],q29=a[3]&b[5],q30=a[3]&b[6],q31=a[3]&b[7],
		q32=a[4]&b[0],q33=a[4]&b[1],q34=a[4]&b[2],q35=a[4]&b[3],q36=a[4]&b[4],q37=a[4]&b[5],q38=a[4]&b[6],q39=a[4]&b[7],
		q40=a[5]&b[0],q41=a[5]&b[1],q42=a[5]&b[2],q43=a[5]&b[3],q44=a[5]&b[4],q45=a[5]&b[5],q46=a[5]&b[6],q47=a[5]&b[7],
		q48=a[6]&b[0],q49=a[6]&b[1],q50=a[6]&b[2],q51=a[6]&b[3],q52=a[6]&b[4],q53=a[6]&b[5],q54=a[6]&b[6],q55=a[6]&b[7],
		q56=a[7]&b[0],q57=a[7]&b[1],q58=a[7]&b[2],q59=a[7]&b[3],q60=a[7]&b[4],q61=a[7]&b[5],q62=a[7]&b[6],q63=a[7]&b[7];


ha x0(q1,q8,p1,c0);
fa x1(q2,q9,q16,s1,c1);
fa x2(q3,q10,q17,s2,c2);
fa x3(q4,q11,q18,s3,c3);
fa x4(q5,q12,q19,s4,c4);
fa x5(q6,q13,q20,s5,c5);
fa x6(q7,q14,q21,s6,c6);


ha x7(s1,c0,p2,c7);
fa x8(q24,s2,c1,s7,c8);
fa x9(q25,s3,c2,s8,c9);
fa x10(q26,s4,c3,s9,c10);
fa x11(q27,s5,c4,s10,c11);
fa x12(q28,s6,c5,s11,c12);
fa x13(q15,q22,c6,s12,c13);

ha x14(s7,c7,p3,c14);
fa x15(q32,s8,c8,s13,c15);
fa x16(q33,s9,c9,s14,c16);
fa x17(q34,s10,c10,s15,c17);
fa x18(q35,s11,c11,s16,c18);
fa x19(q29,s12,c12,s17,c19);
fa x20(q30,q23,c13,s18,c20);

ha x21(s13,c14,p4,c21);
fa x22(q40,s14,c15,s19,c22);
fa x23(q41,s15,c16,s20,c23);
fa x24(q42,s16,c17,s21,c24);
fa x25(q36,s17,c18,s22,c25);
fa x26(q37,s18,c19,s23,c26);
fa x27(q38,q31,c20,s24,c27);

ha x28(s19,c21,p5,c28);
fa x29(q48,s20,c22,s25,c29);
fa x30(q49,s21,c23,s26,c30);
fa x31(q43,s22,c24,s27,c31);
fa x32(q44,s23,c25,s28,c32);
fa x33(q45,s24,c26,s29,c33);
fa x34(q46,q39,c27,s30,c34);

ha x35(s25,c28,p6,c35);
fa x36(q56,s26,c29,s31,c36);
fa x37(q50,s27,c30,s32,c37);
fa x38(q51,s28,c31,s33,c38);
fa x39(q52,s29,c32,s34,c39);
fa x40(q53,s30,c33,s35,c40);
fa x41(q54,q47,c34,s36,c41);

ha x42(s31,c35,p7,c42);
fa x43(q57,s32,c36,s37,c43);
fa x44(q58,s33,c37,s38,c44);
fa x45(q59,s34,c38,s39,c45);
fa x46(q60,s35,c39,s40,c46);
fa x47(q61,s36,c40,s41,c47);
fa x48(q62,q55,c41,s42,c48);

ha x49(s37,c42,p8,c49);
fa x50(s38,c43,c49,p9,c50);
fa x51(s39,c44,c50,p10,c51);
fa x52(s40,c45,c51,p11,c52);
fa x53(s41,c46,c52,p12,c53);
fa x54(s42,c47,c53,p13,c54);
fa x55(q63,c48,c54,p14,p15);

assign out={p15,p14,p13,p12,p11,p10,p9,p8,p7,p6,p5,p4,p3,p2,p1,p0};

endmodule
